import rv32i_types::*;

module ID_EX(
    input clk,
    input rst,
    input load,

    input rv32i_control_word control_word_in,

    input logic [31:0] alu_in,
    input logic [31:0] mdr_in,
    input logic br_en_in,
    input packed_imm imm_in,

    output logic write_en,
    output logic rd,
    output logic [31:0] pc,
    output rv32i_opcode opcode,
    output logic [31:0] alu_out,
    output logic [31:0] mdr_out,
    output logic br_en_out,
    output [31:0] u_imm
);

rv32i_control_word control_word;
logic [31:0] alu, mdr;
logic br_en;
packed_imm imm;

assign rd = control_word.rd;
assign write_en = control_word.write_en;
assign opcode = control_word.opcode;
assign mdr_out = mdr;
assign br_en_out = br_en;
assign u_imm = imm.u_imm;

assign mem_read = control_word.mem_read;
assign mem_write = control_word.mem_write;
assign mem_byte_enable = control_word.mem_byte_enable;

always_ff @(posedge clk)
begin
    if (rst)
    begin
        alu <= 0;
        mdr <= 0;
        br_en <= 0;

        imm.i_imm <= 32'b0;
        imm.s_imm <= 32'b0;
        imm.b_imm <= 32'b0;
        imm.u_imm <= 32'b0;
        imm.j_imm <= 32'b0;

        control_word.opcode <= 0;
        control_word.aluop <= 0;
        control_word.mem_read <= 0;
        control_word.mem_write <= 0;
        control_word.regfilemux_sel <= 0;
        control_word.pcmux_sel <= 0;
        control_word.alumux1_sel <= 0;
        control_word.alumux2_sel <= 0;
        control_word.cmpmux_sel <= 0;
        control_word.rmask <= 0;
        control_word.wmask <= 0;
        control_word.mem_byte_enable <= 0;
        control_word.mem_addr_bits <= 0;
        control_word.rd <= 0;
        control_word.funct3 <= 0;
        control_word.funct7 <= 0;
        control_word.pc <= 0;
    end
    else if (load == 1)
    begin
        control_word <= control_word_in;
        alu <= alu_in;
        mdr <= mdr_in;
        br_en <= br_en_in;
        imm <= imm_in;
    end
    else
    begin
        control_word <= control_word;
        alu <= alu;
        mdr <= mdr;
        br_en <= br_en;
        imm <= imm;
    end
end

endmodule